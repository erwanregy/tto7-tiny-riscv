`ifndef ALU_OPERATIONS_SVH
`define ALU_OPERATIONS_SVH

typedef enum {
    Add,
    Subtract,
    Shift_Left_Logical,
    Set_Less_Than,
    Set_Less_Than_Unsigned,
    Xor,
    Shift_Right_Logical,
    Shift_Right_Arithmetic,
    Or,
    And,
    Invalid
} alu_operation_t;

`endif
