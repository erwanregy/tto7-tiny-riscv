`ifndef OPCODES_SVH
`define OPCODES_SVH

typedef enum logic [6:0] {
    Load_Upper_Immediate = 7'b0110111,
    Add_Upper_Immediate_To_Program_Counter = 7'b0010111,
    Jump_And_Link = 7'b1101111,
    Jump_And_Link_Register = 7'b1100111,
    Branch = 7'b1100011,
    Memory_Access = 7'b0?00011,
    Load = 7'b0000011,
    Store = 7'b0100011,
    Arithmetic = 7'b0?10011,
    Immediate_Arithmetic = 7'b0010011,
    Register_Arithmetic = 7'b0110011,
    Fence = 7'b0001111,
    System = 7'b1110011
} opcode_t;

typedef enum logic [31:0] {
    lui      = 32'b????????????????????____?????_0110111,
    auipc    = 32'b????????????????????____?????_0010111,
    jal      = 32'b????????????????????____?????_1101111,
    jalr     = 32'b????????????__?????_000_?????_1100111,
    beq      = 32'b???????_?????_?????_000_?????_1100011,
    bne      = 32'b???????_?????_?????_001_?????_1100011,
    blt      = 32'b???????_?????_?????_100_?????_1100011,
    bge      = 32'b???????_?????_?????_101_?????_1100011,
    bltu     = 32'b???????_?????_?????_110_?????_1100011,
    bgeu     = 32'b???????_?????_?????_111_?????_1100011,
    lb       = 32'b????????????__?????_000_?????_0000011,
    lh       = 32'b????????????__?????_001_?????_0000011,
    lw       = 32'b????????????__?????_010_?????_0000011,
    lbu      = 32'b????????????__?????_100_?????_0000011,
    lhu      = 32'b????????????__?????_101_?????_0000011,
    sb       = 32'b???????_?????_?????_000_?????_0100011,
    sh       = 32'b???????_?????_?????_001_?????_0100011,
    sw       = 32'b???????_?????_?????_010_?????_0100011,
    addi     = 32'b????????????__?????_000_?????_0010011,
    slti     = 32'b????????????__?????_010_?????_0010011,
    sltiu    = 32'b????????????__?????_011_?????_0010011,
    xori     = 32'b????????????__?????_100_?????_0010011,
    ori      = 32'b????????????__?????_110_?????_0010011,
    andi     = 32'b????????????__?????_111_?????_0010011,
    slli     = 32'b0000000_?????_?????_001_?????_0010011,
    srli     = 32'b0000000_?????_?????_101_?????_0010011,
    srai     = 32'b0100000_?????_?????_101_?????_0010011,
    add      = 32'b0000000_?????_?????_000_?????_0110011,
    sub      = 32'b0100000_?????_?????_000_?????_0110011,
    sll      = 32'b0000000_?????_?????_001_?????_0110011,
    slt      = 32'b0000000_?????_?????_010_?????_0110011,
    sltu     = 32'b0000000_?????_?????_011_?????_0110011,
    xor_     = 32'b0000000_?????_?????_100_?????_0110011,
    srl      = 32'b0000000_?????_?????_101_?????_0110011,
    sra      = 32'b0100000_?????_?????_101_?????_0110011,
    or_      = 32'b0000000_?????_?????_110_?????_0110011,
    and_     = 32'b0000000_?????_?????_111_?????_0110011,
    fence    = 32'b0000000_?????_?????_000_?????_0001111,
    fence_i  = 32'b0000000_?????_?????_001_?????_0001111,
    ecall    = 32'b000000000000__00000_000_00000_1110011,
    ebreak   = 32'b000000000001__00000_000_00000_1110011,
    csrrw    = 32'b?????????????????___001_?????_1110011,
    csrrs    = 32'b?????????????????___010_?????_1110011,
    csrrc    = 32'b?????????????????___011_?????_1110011,
    csrrwi   = 32'b?????????????????___101_?????_1110011,
    csrrsi   = 32'b?????????????????___110_?????_1110011,
    csrrci   = 32'b?????????????????___111_?????_1110011,
    nop      = 32'b?????????????????????????_____0000000,
    invalid  = 0
} operation_t;

`endif
